module add_sub;

  reg [4:0] a_1, a_2, b_2, a_3, b_3;
  reg [1:0] b_2;
  reg [31:0] 
  
