`include "struct_types.sv"
import float_struct::*;


module shift_reg_for_struct(
  input               clk,
  input               rst,

);





endmodule
