module division();



endmodule
