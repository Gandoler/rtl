module division_test();



endmodule
