module mul



endmodule
