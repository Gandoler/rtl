package float_types_pkg;
typedef struct packed {
  logic        sign;
  logic [7:0]  exp;
  logic [23:0] mant;
} float_point_num;

typedef enum logic [1:0]{
  OK_state         = 2'b00,
  NAN_or_INF = 2'b01,
  ZERO_res = 2'b10
} num_status;
endpackage
