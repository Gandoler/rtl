module mul();

logic [7:0] mul1 ,mul2;

assign mul1 = 3'd7 * 5'd20;
assign mul2 = 3'd7 * 5'd31;

endmodule
