module div_block(
  input logic R,
  input logic B,
  input logic C_in,

  output logic C_out,
  output logic D,
  output logic B_out,
  output logic R_out
);
