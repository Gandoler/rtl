module FDCE(
    input  logic C,
    input  logic CE,
    input  logic PRE,
    input  logic D,
    output logic Q
);




endmodule
